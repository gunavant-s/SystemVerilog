module add(add_if inf);
  
  assign inf.sum = inf.a | inf.b; //Here we are not declaring variables
  
endmodule
